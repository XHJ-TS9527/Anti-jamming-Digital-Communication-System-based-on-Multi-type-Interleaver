library ieee;
use ieee.std_logic_1164.all;
entity circle_address_selector is
	port(guide:in std_logic_vector(7 downto 0);
		 CS:in std_logic; --chip select signal
		 W_address:out std_logic_vector(7 downto 0));
end circle_address_selector;
architecture dataflow of circle_address_selector is
signal WR_add:std_logic_vector(7 downto 0);
begin
	W_address<=WR_add when (CS='1') else (others=>'Z');
	with guide select
		WR_add<="00000000" when "00000000",
				"00010001" when "00000001",
				"00100010" when "00000010",
				"00110011" when "00000011",
				"01000100" when "00000100",
				"01010101" when "00000101",
				"01100110" when "00000110",
				"01110111" when "00000111",
				"10001000" when "00001000",
				"10011001" when "00001001",
				"10101010" when "00001010",
				"10111011" when "00001011",
				"10111100" when "00001100",
				"10111101" when "00001101",
				"10111110" when "00001110",
				"10111111" when "00001111",
				"11000000" when "00010000",
				"11000001" when "00010001",
				"11000010" when "00010010",
				"11000011" when "00010011",
				"11000100" when "00010100",
				"11000101" when "00010101",
				"11000110" when "00010110",
				"11000111" when "00010111",
				"11001000" when "00011000",
				"11001001" when "00011001",
				"11001010" when "00011010",
				"11001011" when "00011011",
				"10111010" when "00011100",
				"10101001" when "00011101",
				"10011000" when "00011110",
				"10000111" when "00011111",
				"01110110" when "00100000",
				"01100101" when "00100001",
				"01010100" when "00100010",
				"01000011" when "00100011",
				"00110010" when "00100100",
				"00100001" when "00100101",
				"00010000" when "00100110",
				"00001111" when "00100111",
				"00001110" when "00101000",
				"00001101" when "00101001",
				"00001100" when "00101010",
				"00001011" when "00101011",
				"00001010" when "00101100",
				"00001001" when "00101101",
				"00001000" when "00101110",
				"00000111" when "00101111",
				"00000110" when "00110000",
				"00000101" when "00110001",
				"00000100" when "00110010",
				"00000011" when "00110011",
				"00000010" when "00110100",
				"00000001" when "00110101",
				"00010010" when "00110110",
				"00100011" when "00110111",
				"00110100" when "00111000",
				"01000101" when "00111001",
				"01010110" when "00111010",
				"01100111" when "00111011",
				"01111000" when "00111100",
				"10001001" when "00111101",
				"10011010" when "00111110",
				"10101011" when "00111111",
				"10101100" when "01000000",
				"10101101" when "01000001",
				"10101110" when "01000010",
				"10101111" when "01000011",
				"10110000" when "01000100",
				"10110001" when "01000101",
				"10110010" when "01000110",
				"10110011" when "01000111",
				"10110100" when "01001000",
				"10110101" when "01001001",
				"10110110" when "01001010",
				"10110111" when "01001011",
				"10111000" when "01001100",
				"10111001" when "01001101",
				"10101000" when "01001110",
				"10010111" when "01001111",
				"10000110" when "01010000",
				"01110101" when "01010001",
				"01100100" when "01010010",
				"01010011" when "01010011",
				"01000010" when "01010100",
				"00110001" when "01010101",
				"00100000" when "01010110",
				"00011111" when "01010111",
				"00011110" when "01011000",
				"00011101" when "01011001",
				"00011100" when "01011010",
				"00011011" when "01011011",
				"00011010" when "01011100",
				"00011001" when "01011101",
				"00011000" when "01011110",
				"00010111" when "01011111",
				"00010110" when "01100000",
				"00010101" when "01100001",
				"00010100" when "01100010",
				"00010011" when "01100011",
				"00100100" when "01100100",
				"00110101" when "01100101",
				"01000110" when "01100110",
				"01010111" when "01100111",
				"01101000" when "01101000",
				"01111001" when "01101001",
				"10001010" when "01101010",
				"10011011" when "01101011",
				"10011100" when "01101100",
				"10011101" when "01101101",
				"10011110" when "01101110",
				"10011111" when "01101111",
				"10100000" when "01110000",
				"10100001" when "01110001",
				"10100010" when "01110010",
				"10100011" when "01110011",
				"10100100" when "01110100",
				"10100101" when "01110101",
				"10100110" when "01110110",
				"10100111" when "01110111",
				"10010110" when "01111000",
				"10000101" when "01111001",
				"01110100" when "01111010",
				"01100011" when "01111011",
				"01010010" when "01111100",
				"01000001" when "01111101",
				"00110000" when "01111110",
				"00101111" when "01111111",
				"00101110" when "10000000",
				"00101101" when "10000001",
				"00101100" when "10000010",
				"00101011" when "10000011",
				"00101010" when "10000100",
				"00101001" when "10000101",
				"00101000" when "10000110",
				"00100111" when "10000111",
				"00100110" when "10001000",
				"00100101" when "10001001",
				"00110110" when "10001010",
				"01000111" when "10001011",
				"01011000" when "10001100",
				"01101001" when "10001101",
				"01111010" when "10001110",
				"10001011" when "10001111",
				"10001100" when "10010000",
				"10001101" when "10010001",
				"10001110" when "10010010",
				"10001111" when "10010011",
				"10010000" when "10010100",
				"10010001" when "10010101",
				"10010010" when "10010110",
				"10010011" when "10010111",
				"10010100" when "10011000",
				"10010101" when "10011001",
				"10000100" when "10011010",
				"01110011" when "10011011",
				"01100010" when "10011100",
				"01010001" when "10011101",
				"01000000" when "10011110",
				"00111111" when "10011111",
				"00111110" when "10100000",
				"00111101" when "10100001",
				"00111100" when "10100010",
				"00111011" when "10100011",
				"00111010" when "10100100",
				"00111001" when "10100101",
				"00111000" when "10100110",
				"00110111" when "10100111",
				"01001000" when "10101000",
				"01011001" when "10101001",
				"01101010" when "10101010",
				"01111011" when "10101011",
				"01111100" when "10101100",
				"01111101" when "10101101",
				"01111110" when "10101110",
				"01111111" when "10101111",
				"10000000" when "10110000",
				"10000001" when "10110001",
				"10000010" when "10110010",
				"10000011" when "10110011",
				"01110010" when "10110100",
				"01100001" when "10110101",
				"01010000" when "10110110",
				"01001111" when "10110111",
				"01001110" when "10111000",
				"01001101" when "10111001",
				"01001100" when "10111010",
				"01001011" when "10111011",
				"01001010" when "10111100",
				"01001001" when "10111101",
				"01011010" when "10111110",
				"01101011" when "10111111",
				"01101100" when "11000000",
				"01101101" when "11000001",
				"01101110" when "11000010",
				"01101111" when "11000011",
				"01110000" when "11000100",
				"01110001" when "11000101",
				"01100000" when "11000110",
				"01011111" when "11000111",
				"01011110" when "11001000",
				"01011101" when "11001001",
				"01011100" when "11001010",
				"01011011" when "11001011",
				"00000000" when others;
end dataflow;