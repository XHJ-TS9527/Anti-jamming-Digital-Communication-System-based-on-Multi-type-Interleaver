library ieee;
use ieee.std_logic_1164.all;
entity oddeven_address_selector is
	port(guide:in std_logic_vector(7 downto 0);
		 CS:in std_logic; --chip select signal
		 W_address:out std_logic_vector(7 downto 0));
end oddeven_address_selector;
architecture dataflow of oddeven_address_selector is
signal WR_add:std_logic_vector(7 downto 0);
begin
	W_address<=WR_add when (CS='1') else (others=>'Z');
	with guide select
		WR_add<="00000000" when "00000000",
				"00000010" when "00000001",
				"00000100" when "00000010",
				"00000110" when "00000011",
				"00001000" when "00000100",
				"00001010" when "00000101",
				"00001100" when "00000110",
				"00001110" when "00000111",
				"00010000" when "00001000",
				"00010010" when "00001001",
				"00010100" when "00001010",
				"00010110" when "00001011",
				"00011000" when "00001100",
				"00011010" when "00001101",
				"00011100" when "00001110",
				"00011110" when "00001111",
				"00100000" when "00010000",
				"00100010" when "00010001",
				"00100100" when "00010010",
				"00100110" when "00010011",
				"00101000" when "00010100",
				"00101010" when "00010101",
				"00101100" when "00010110",
				"00101110" when "00010111",
				"00110000" when "00011000",
				"00110010" when "00011001",
				"00110100" when "00011010",
				"00110110" when "00011011",
				"00111000" when "00011100",
				"00111010" when "00011101",
				"00111100" when "00011110",
				"00111110" when "00011111",
				"01000000" when "00100000",
				"01000010" when "00100001",
				"01000100" when "00100010",
				"01000110" when "00100011",
				"01001000" when "00100100",
				"01001010" when "00100101",
				"01001100" when "00100110",
				"01001110" when "00100111",
				"01010000" when "00101000",
				"01010010" when "00101001",
				"01010100" when "00101010",
				"01010110" when "00101011",
				"01011000" when "00101100",
				"01011010" when "00101101",
				"01011100" when "00101110",
				"01011110" when "00101111",
				"01100000" when "00110000",
				"01100010" when "00110001",
				"01100100" when "00110010",
				"01100110" when "00110011",
				"01101000" when "00110100",
				"01101010" when "00110101",
				"01101100" when "00110110",
				"01101110" when "00110111",
				"01110000" when "00111000",
				"01110010" when "00111001",
				"01110100" when "00111010",
				"01110110" when "00111011",
				"01111000" when "00111100",
				"01111010" when "00111101",
				"01111100" when "00111110",
				"01111110" when "00111111",
				"10000000" when "01000000",
				"10000010" when "01000001",
				"10000100" when "01000010",
				"10000110" when "01000011",
				"10001000" when "01000100",
				"10001010" when "01000101",
				"10001100" when "01000110",
				"10001110" when "01000111",
				"10010000" when "01001000",
				"10010010" when "01001001",
				"10010100" when "01001010",
				"10010110" when "01001011",
				"10011000" when "01001100",
				"10011010" when "01001101",
				"10011100" when "01001110",
				"10011110" when "01001111",
				"10100000" when "01010000",
				"10100010" when "01010001",
				"10100100" when "01010010",
				"10100110" when "01010011",
				"10101000" when "01010100",
				"10101010" when "01010101",
				"10101100" when "01010110",
				"10101110" when "01010111",
				"10110000" when "01011000",
				"10110010" when "01011001",
				"10110100" when "01011010",
				"10110110" when "01011011",
				"10111000" when "01011100",
				"10111010" when "01011101",
				"10111100" when "01011110",
				"10111110" when "01011111",
				"11000000" when "01100000",
				"11000010" when "01100001",
				"11000100" when "01100010",
				"11000110" when "01100011",
				"11001000" when "01100100",
				"11001010" when "01100101",
				"00000001" when "01100110",
				"00000011" when "01100111",
				"00000101" when "01101000",
				"00000111" when "01101001",
				"00001001" when "01101010",
				"00001011" when "01101011",
				"00001101" when "01101100",
				"00001111" when "01101101",
				"00010001" when "01101110",
				"00010011" when "01101111",
				"00010101" when "01110000",
				"00010111" when "01110001",
				"00011001" when "01110010",
				"00011011" when "01110011",
				"00011101" when "01110100",
				"00011111" when "01110101",
				"00100001" when "01110110",
				"00100011" when "01110111",
				"00100101" when "01111000",
				"00100111" when "01111001",
				"00101001" when "01111010",
				"00101011" when "01111011",
				"00101101" when "01111100",
				"00101111" when "01111101",
				"00110001" when "01111110",
				"00110011" when "01111111",
				"00110101" when "10000000",
				"00110111" when "10000001",
				"00111001" when "10000010",
				"00111011" when "10000011",
				"00111101" when "10000100",
				"00111111" when "10000101",
				"01000001" when "10000110",
				"01000011" when "10000111",
				"01000101" when "10001000",
				"01000111" when "10001001",
				"01001001" when "10001010",
				"01001011" when "10001011",
				"01001101" when "10001100",
				"01001111" when "10001101",
				"01010001" when "10001110",
				"01010011" when "10001111",
				"01010101" when "10010000",
				"01010111" when "10010001",
				"01011001" when "10010010",
				"01011011" when "10010011",
				"01011101" when "10010100",
				"01011111" when "10010101",
				"01100001" when "10010110",
				"01100011" when "10010111",
				"01100101" when "10011000",
				"01100111" when "10011001",
				"01101001" when "10011010",
				"01101011" when "10011011",
				"01101101" when "10011100",
				"01101111" when "10011101",
				"01110001" when "10011110",
				"01110011" when "10011111",
				"01110101" when "10100000",
				"01110111" when "10100001",
				"01111001" when "10100010",
				"01111011" when "10100011",
				"01111101" when "10100100",
				"01111111" when "10100101",
				"10000001" when "10100110",
				"10000011" when "10100111",
				"10000101" when "10101000",
				"10000111" when "10101001",
				"10001001" when "10101010",
				"10001011" when "10101011",
				"10001101" when "10101100",
				"10001111" when "10101101",
				"10010001" when "10101110",
				"10010011" when "10101111",
				"10010101" when "10110000",
				"10010111" when "10110001",
				"10011001" when "10110010",
				"10011011" when "10110011",
				"10011101" when "10110100",
				"10011111" when "10110101",
				"10100001" when "10110110",
				"10100011" when "10110111",
				"10100101" when "10111000",
				"10100111" when "10111001",
				"10101001" when "10111010",
				"10101011" when "10111011",
				"10101101" when "10111100",
				"10101111" when "10111101",
				"10110001" when "10111110",
				"10110011" when "10111111",
				"10110101" when "11000000",
				"10110111" when "11000001",
				"10111001" when "11000010",
				"10111011" when "11000011",
				"10111101" when "11000100",
				"10111111" when "11000101",
				"11000001" when "11000110",
				"11000011" when "11000111",
				"11000101" when "11001000",
				"11000111" when "11001001",
				"11001001" when "11001010",
				"11001011" when "11001011",
				"00000000" when others;
end dataflow;