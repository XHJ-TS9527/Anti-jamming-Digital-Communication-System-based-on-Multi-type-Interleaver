library ieee;
use ieee.std_logic_1164.all;
entity interdigital_address_selector is
	port(guide:in std_logic_vector(7 downto 0);
		 CS:in std_logic; --chip select signal
		 W_address:out std_logic_vector(7 downto 0));
end interdigital_address_selector;
architecture dataflow of interdigital_address_selector is
signal WR_add:std_logic_vector(7 downto 0);
begin
	W_address<=WR_add when (CS='1') else (others=>'Z');
	with guide select
		WR_add<="00000000" when "00000000",
				"00010001" when "00000001",
				"00100010" when "00000010",
				"00110011" when "00000011",
				"01000100" when "00000100",
				"01010101" when "00000101",
				"01100110" when "00000110",
				"01110111" when "00000111",
				"10001000" when "00001000",
				"10011001" when "00001001",
				"10101010" when "00001010",
				"10111011" when "00001011",
				"10111100" when "00001100",
				"10101011" when "00001101",
				"10011010" when "00001110",
				"10001001" when "00001111",
				"01111000" when "00010000",
				"01100111" when "00010001",
				"01010110" when "00010010",
				"01000101" when "00010011",
				"00110100" when "00010100",
				"00100011" when "00010101",
				"00010010" when "00010110",
				"00000001" when "00010111",
				"00000010" when "00011000",
				"00010011" when "00011001",
				"00100100" when "00011010",
				"00110101" when "00011011",
				"01000110" when "00011100",
				"01010111" when "00011101",
				"01101000" when "00011110",
				"01111001" when "00011111",
				"10001010" when "00100000",
				"10011011" when "00100001",
				"10101100" when "00100010",
				"10111101" when "00100011",
				"10111110" when "00100100",
				"10101101" when "00100101",
				"10011100" when "00100110",
				"10001011" when "00100111",
				"01111010" when "00101000",
				"01101001" when "00101001",
				"01011000" when "00101010",
				"01000111" when "00101011",
				"00110110" when "00101100",
				"00100101" when "00101101",
				"00010100" when "00101110",
				"00000011" when "00101111",
				"00000100" when "00110000",
				"00010101" when "00110001",
				"00100110" when "00110010",
				"00110111" when "00110011",
				"01001000" when "00110100",
				"01011001" when "00110101",
				"01101010" when "00110110",
				"01111011" when "00110111",
				"10001100" when "00111000",
				"10011101" when "00111001",
				"10101110" when "00111010",
				"10111111" when "00111011",
				"11000000" when "00111100",
				"10101111" when "00111101",
				"10011110" when "00111110",
				"10001101" when "00111111",
				"01111100" when "01000000",
				"01101011" when "01000001",
				"01011010" when "01000010",
				"01001001" when "01000011",
				"00111000" when "01000100",
				"00100111" when "01000101",
				"00010110" when "01000110",
				"00000101" when "01000111",
				"00000110" when "01001000",
				"00010111" when "01001001",
				"00101000" when "01001010",
				"00111001" when "01001011",
				"01001010" when "01001100",
				"01011011" when "01001101",
				"01101100" when "01001110",
				"01111101" when "01001111",
				"10001110" when "01010000",
				"10011111" when "01010001",
				"10110000" when "01010010",
				"11000001" when "01010011",
				"11000010" when "01010100",
				"10110001" when "01010101",
				"10100000" when "01010110",
				"10001111" when "01010111",
				"01111110" when "01011000",
				"01101101" when "01011001",
				"01011100" when "01011010",
				"01001011" when "01011011",
				"00111010" when "01011100",
				"00101001" when "01011101",
				"00011000" when "01011110",
				"00000111" when "01011111",
				"00001000" when "01100000",
				"00011001" when "01100001",
				"00101010" when "01100010",
				"00111011" when "01100011",
				"01001100" when "01100100",
				"01011101" when "01100101",
				"01101110" when "01100110",
				"01111111" when "01100111",
				"10010000" when "01101000",
				"10100001" when "01101001",
				"10110010" when "01101010",
				"11000011" when "01101011",
				"11000100" when "01101100",
				"10110011" when "01101101",
				"10100010" when "01101110",
				"10010001" when "01101111",
				"10000000" when "01110000",
				"01101111" when "01110001",
				"01011110" when "01110010",
				"01001101" when "01110011",
				"00111100" when "01110100",
				"00101011" when "01110101",
				"00011010" when "01110110",
				"00001001" when "01110111",
				"00001010" when "01111000",
				"00011011" when "01111001",
				"00101100" when "01111010",
				"00111101" when "01111011",
				"01001110" when "01111100",
				"01011111" when "01111101",
				"01110000" when "01111110",
				"10000001" when "01111111",
				"10010010" when "10000000",
				"10100011" when "10000001",
				"10110100" when "10000010",
				"11000101" when "10000011",
				"11000110" when "10000100",
				"10110101" when "10000101",
				"10100100" when "10000110",
				"10010011" when "10000111",
				"10000010" when "10001000",
				"01110001" when "10001001",
				"01100000" when "10001010",
				"01001111" when "10001011",
				"00111110" when "10001100",
				"00101101" when "10001101",
				"00011100" when "10001110",
				"00001011" when "10001111",
				"00001100" when "10010000",
				"00011101" when "10010001",
				"00101110" when "10010010",
				"00111111" when "10010011",
				"01010000" when "10010100",
				"01100001" when "10010101",
				"01110010" when "10010110",
				"10000011" when "10010111",
				"10010100" when "10011000",
				"10100101" when "10011001",
				"10110110" when "10011010",
				"11000111" when "10011011",
				"11001000" when "10011100",
				"10110111" when "10011101",
				"10100110" when "10011110",
				"10010101" when "10011111",
				"10000100" when "10100000",
				"01110011" when "10100001",
				"01100010" when "10100010",
				"01010001" when "10100011",
				"01000000" when "10100100",
				"00101111" when "10100101",
				"00011110" when "10100110",
				"00001101" when "10100111",
				"00001110" when "10101000",
				"00011111" when "10101001",
				"00110000" when "10101010",
				"01000001" when "10101011",
				"01010010" when "10101100",
				"01100011" when "10101101",
				"01110100" when "10101110",
				"10000101" when "10101111",
				"10010110" when "10110000",
				"10100111" when "10110001",
				"10111000" when "10110010",
				"11001001" when "10110011",
				"11001010" when "10110100",
				"10111001" when "10110101",
				"10101000" when "10110110",
				"10010111" when "10110111",
				"10000110" when "10111000",
				"01110101" when "10111001",
				"01100100" when "10111010",
				"01010011" when "10111011",
				"01000010" when "10111100",
				"00110001" when "10111101",
				"00100000" when "10111110",
				"00001111" when "10111111",
				"00010000" when "11000000",
				"00100001" when "11000001",
				"00110010" when "11000010",
				"01000011" when "11000011",
				"01010100" when "11000100",
				"01100101" when "11000101",
				"01110110" when "11000110",
				"10000111" when "11000111",
				"10011000" when "11001000",
				"10101001" when "11001001",
				"10111010" when "11001010",
				"11001011" when "11001011",
				"00000000" when others;
end dataflow;