library ieee;
use ieee.std_logic_1164.all;
entity pseudorandom_address_selector is
	port(guide:in std_logic_vector(7 downto 0);
		 CS:in std_logic; --chip select signal
		 W_address:out std_logic_vector(7 downto 0));
end pseudorandom_address_selector;
architecture dataflow of pseudorandom_address_selector is
signal WR_add:std_logic_vector(7 downto 0);
begin
	W_address<=WR_add when (CS='1') else (others=>'Z');
	with guide select
		WR_add<="01110110" when "00000000",
				"01011110" when "00000001",
				"10101001" when "00000010",
				"00011011" when "00000011",
				"00100011" when "00000100",
				"00010001" when "00000101",
				"10101010" when "00000110",
				"00011101" when "00000111",
				"10010011" when "00001000",
				"01010111" when "00001001",
				"10100101" when "00001010",
				"01010110" when "00001011",
				"10001101" when "00001100",
				"01110010" when "00001101",
				"10111001" when "00001110",
				"01101011" when "00001111",
				"01111010" when "00010000",
				"10100000" when "00010001",
				"00011110" when "00010010",
				"00000001" when "00010011",
				"01110100" when "00010100",
				"10011011" when "00010101",
				"00110010" when "00010110",
				"10001111" when "00010111",
				"01011011" when "00011000",
				"10100001" when "00011001",
				"10000011" when "00011010",
				"00111111" when "00011011",
				"00001011" when "00011100",
				"10000111" when "00011101",
				"10000010" when "00011110",
				"01000000" when "00011111",
				"01101110" when "00100000",
				"00000110" when "00100001",
				"01100000" when "00100010",
				"00110001" when "00100011",
				"01100100" when "00100100",
				"10101011" when "00100101",
				"00011001" when "00100110",
				"10000000" when "00100111",
				"10110101" when "00101000",
				"10010000" when "00101001",
				"00101000" when "00101010",
				"10110011" when "00101011",
				"01001000" when "00101100",
				"00110111" when "00101101",
				"01101100" when "00101110",
				"10100110" when "00101111",
				"10001110" when "00110000",
				"10010001" when "00110001",
				"10011110" when "00110010",
				"01000101" when "00110011",
				"01001001" when "00110100",
				"01000011" when "00110101",
				"00111001" when "00110110",
				"01000001" when "00110111",
				"01111100" when "00111000",
				"01100110" when "00111001",
				"10000001" when "00111010",
				"00101110" when "00111011",
				"00011100" when "00111100",
				"00000010" when "00111101",
				"01010001" when "00111110",
				"10110001" when "00111111",
				"10111111" when "01000000",
				"01100010" when "01000001",
				"00100001" when "01000010",
				"01011111" when "01000011",
				"10011000" when "01000100",
				"00110101" when "01000101",
				"01000111" when "01000110",
				"11001000" when "01000111",
				"10001010" when "01001000",
				"01001100" when "01001001",
				"10100111" when "01001010",
				"10110110" when "01001011",
				"10011010" when "01001100",
				"11000101" when "01001101",
				"01010100" when "01001110",
				"00100101" when "01001111",
				"10011101" when "01010000",
				"00010111" when "01010001",
				"01111011" when "01010010",
				"10001100" when "01010011",
				"10011111" when "01010100",
				"10010010" when "01010101",
				"00001100" when "01010110",
				"01111110" when "01010111",
				"10111101" when "01011000",
				"00100100" when "01011001",
				"01110011" when "01011010",
				"00101010" when "01011011",
				"10111110" when "01011100",
				"01101010" when "01011101",
				"10101111" when "01011110",
				"01011101" when "01011111",
				"01001011" when "01100000",
				"00001001" when "01100001",
				"10111100" when "01100010",
				"10010111" when "01100011",
				"00101001" when "01100100",
				"10010110" when "01100101",
				"00110011" when "01100110",
				"00111010" when "01100111",
				"11000000" when "01101000",
				"11000001" when "01101001",
				"10001011" when "01101010",
				"01100011" when "01101011",
				"01011000" when "01101100",
				"11000111" when "01101101",
				"01110000" when "01101110",
				"00000011" when "01101111",
				"10110000" when "01110000",
				"00111110" when "01110001",
				"01001111" when "01110010",
				"10000110" when "01110011",
				"11001011" when "01110100",
				"01010101" when "01110101",
				"01011100" when "01110110",
				"10100100" when "01110111",
				"10000101" when "01111000",
				"01001110" when "01111001",
				"00110110" when "01111010",
				"01100101" when "01111011",
				"01001010" when "01111100",
				"10001001" when "01111101",
				"10110111" when "01111110",
				"00000000" when "01111111",
				"11000100" when "10000000",
				"00101011" when "10000001",
				"10101110" when "10000010",
				"10101100" when "10000011",
				"01100111" when "10000100",
				"00110000" when "10000101",
				"00011000" when "10000110",
				"00010000" when "10000111",
				"00010100" when "10001000",
				"00101111" when "10001001",
				"10110100" when "10001010",
				"01101000" when "10001011",
				"00100000" when "10001100",
				"00111011" when "10001101",
				"00011010" when "10001110",
				"00101100" when "10001111",
				"10101101" when "10010000",
				"00010110" when "10010001",
				"10110010" when "10010010",
				"01101001" when "10010011",
				"00111000" when "10010100",
				"01010011" when "10010101",
				"00101101" when "10010110",
				"01010010" when "10010111",
				"00010101" when "10011000",
				"00100110" when "10011001",
				"01110111" when "10011010",
				"10111011" when "10011011",
				"01011001" when "10011100",
				"10111000" when "10011101",
				"10011100" when "10011110",
				"00001110" when "10011111",
				"01100001" when "10100000",
				"11000011" when "10100001",
				"00100111" when "10100010",
				"01111101" when "10100011",
				"00001010" when "10100100",
				"11000110" when "10100101",
				"01000100" when "10100110",
				"01111000" when "10100111",
				"11000010" when "10101000",
				"10101000" when "10101001",
				"00011111" when "10101010",
				"01101111" when "10101011",
				"01001101" when "10101100",
				"01000010" when "10101101",
				"00010010" when "10101110",
				"10001000" when "10101111",
				"01111001" when "10110000",
				"10000100" when "10110001",
				"11001010" when "10110010",
				"00111100" when "10110011",
				"10011001" when "10110100",
				"10010100" when "10110101",
				"01111111" when "10110110",
				"01101101" when "10110111",
				"00001101" when "10111000",
				"01010000" when "10111001",
				"01000110" when "10111010",
				"10111010" when "10111011",
				"00010011" when "10111100",
				"01011010" when "10111101",
				"11001001" when "10111110",
				"10100010" when "10111111",
				"10010101" when "11000000",
				"00100010" when "11000001",
				"10100011" when "11000010",
				"00001000" when "11000011",
				"00000100" when "11000100",
				"00111101" when "11000101",
				"00001111" when "11000110",
				"00110100" when "11000111",
				"01110101" when "11001000",
				"00000101" when "11001001",
				"00000111" when "11001010",
				"01110001" when "11001011",
				"01110110" when others;
end dataflow;